`timescale 1ns / 1ps

module tcp_top(
    input                               clk                        ,
    input                               rst_n                      
);
                                                                   
                                                                   
endmodule